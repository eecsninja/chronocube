// Copyright (C) 2013 Simon Que
//
// This file is part of ChronoCube.
//
// ChronoCube is free software: you can redistribute it and/or modify
// it under the terms of the GNU Lesser General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// ChronoCube is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public License
// along with ChronoCube.  If not, see <http://www.gnu.org/licenses/>.


// Top-level ChronoCube module.

`include "registers.vh"
`include "tile_registers.vh"

`define MPU_ADDR_WIDTH 16
`define MPU_DATA_WIDTH 16

`define VRAM_ADDR_WIDTH 16
`define VRAM_DATA_WIDTH 16

`define RGB_COLOR_DEPTH 18

`define DISPLAY_HCOUNT_WIDTH 10
`define DISPLAY_VCOUNT_WIDTH 10

`define PAL_ADDR_BASE   'h0800
`define PAL_ADDR_LENGTH    512

`define PAL_ADDR_WIDTH 10
`define PAL_DATA_WIDTH 24
`define MPU_DATA_WIDTH 16
`define NUM_PAL_CHANNELS 3

module ChronoCube(clk, _reset, _int,
                  _mpu_rd, _mpu_wr, _mpu_en, _mpu_be, mpu_addr, mpu_data,
                  _vram_en, _vram_rd, _vram_wr, _vram_be, vram_addr, vram_data,
                  vga_vsync, vga_hsync, vga_rgb);

  input clk;                // System clock

  input _reset;             // Reset (active low)
  input _int;               // Interrupt (active low)

  // MPU-side interface
  input _mpu_en;            // Enable access (active low)
  input _mpu_rd;            // Read enable (active low)
  input _mpu_wr;            // Write enable (active low)
  input [1:0] _mpu_be;      // Byte enable (active low)
  input [`MPU_ADDR_WIDTH-1:0] mpu_addr;  // Address bus
  inout [`MPU_DATA_WIDTH-1:0] mpu_data;  // Data bus

  // VRAM interface
  output _vram_en;          // Enable access (active low)
  output _vram_rd;          // Read enable (active low)
  output _vram_wr;          // Write enable (active low)
  output [1:0] _vram_be;    // Byte enable (active low)
  output [`VRAM_ADDR_WIDTH-1:0] vram_addr;   // Address bus
  inout [`VRAM_DATA_WIDTH-1:0]  vram_data;   // Data bus

  // VGA display interface
  // Note that Hsync and Vsync are active low for some modes and active high for
  // others.
  output vga_vsync;        // Hsync
  output vga_hsync;        // Vsync
  output [`RGB_COLOR_DEPTH-1:0] vga_rgb;   // RGB data

  // VGA signal generator
  // Counters for the position of the refresh.
  wire [`DISPLAY_HCOUNT_WIDTH-1:0] h_pos;
  wire [`DISPLAY_VCOUNT_WIDTH-1:0] v_pos;
  // Signals to indicate that refresh is in an off-screen area.
  wire hblank;
  wire vblank;
  DisplayController #(.HCOUNT_WIDTH(`DISPLAY_HCOUNT_WIDTH),
                      .VCOUNT_WIDTH(`DISPLAY_VCOUNT_WIDTH))
      display(.clk(clk),
              ._reset(_reset),
              .v_pos(v_pos),
              .h_pos(h_pos),
              .hsync(vga_hsync),
              .vsync(vga_vsync),
              .vblank(vblank),
              .hblank(hblank));

  // Graphics processor
  // TODO: add switching between 16-bit full color and 8-bit palettes.
  wire [`VRAM_ADDR_WIDTH-1:0] ren_bus_addr;
  wire [`VRAM_DATA_WIDTH-1:0] ren_bus_data;
  wire _ren_bus_en;
  wire _ren_bus_rd;
  wire _ren_bus_wr;
  wire [1:0] _ren_bus_be;
  wire [`RGB_COLOR_DEPTH-1:0] ren_rgb_out;

  wire [`MPU_DATA_WIDTH-1:0] pal_data_out;
  wire [`MPU_DATA_WIDTH-1:0] reg_data_out;
  assign mpu_data = (_mpu_rd | _mpu_en) ? {`MPU_DATA_WIDTH {1'bz}} :
                    (palette_select  ? pal_data_out :
                    (map_select      ? map_data_out :
                    (main_reg_select ? reg_data_out :
                    {`MPU_DATA_WIDTH {1'b0}})));

  // Palette interface
  wire palette_select = (mpu_addr >= `PAL_ADDR_BASE) &
                        (mpu_addr < `PAL_ADDR_BASE + `PAL_ADDR_LENGTH);
  wire pal_wr = palette_select & ~_mpu_wr;
  wire pal_rd = palette_select & ~_mpu_rd;

  wire [`NUM_PAL_CHANNELS-1:0] pal_byte_en;
  assign pal_byte_en[0] = (mpu_addr[0] == 0) & ~_mpu_be[0];
  assign pal_byte_en[1] = (mpu_addr[0] == 0) & ~_mpu_be[1];
  assign pal_byte_en[2] = (mpu_addr[0] == 1) & ~_mpu_be[0];

  wire [`NUM_PAL_CHANNELS*8-1:0] pal_data_out_temp;
  assign pal_data_out = (mpu_addr[0] == 0) ? pal_data_out_temp[15:0]
                                           : pal_data_out_temp[23:16];

  wire [`PAL_ADDR_WIDTH-1:0] ren_pal_addr;
  wire [`NUM_PAL_CHANNELS*8-1:0] ren_pal_data_out;
  Palette #(.NUM_CHANNELS(`NUM_PAL_CHANNELS)) palette(
      .clk_a(clk),
      .wr_a(pal_wr),
      .rd_a(pal_rd),
      .addr_a(mpu_addr >> 1),
      .data_in_a({mpu_data, mpu_data}),
      .data_out_a(pal_data_out_temp),
      .byte_en_a(pal_byte_en),
      .clk_b(clk),
      .wr_b(0),
      .rd_b(1),
      .addr_b(ren_pal_addr),
      .data_out_b(ren_pal_data_out)
      );

  // Tile map
  wire map_select = (mpu_addr >= `TILEMAP_ADDR_BASE) &
                    (mpu_addr < `TILEMAP_ADDR_BASE + `TILEMAP_ADDR_LENGTH);
  wire map_wr = map_select & ~_mpu_wr;
  wire map_rd = map_select & ~_mpu_rd;
  wire [1:0] map_be = ~_mpu_be;
  wire [`MPU_DATA_WIDTH-1:0] map_data_out;
  tilemap_ram_4Kx16 tilemap(
      .clock_a(clk),
      .clock_b(clk),
      .address_a(mpu_addr),
      .byteena_a(map_be),
      .data_a(mpu_data),
      .data_b(0),
      .rden_a(map_rd),
      .rden_b(0),
      .wren_a(map_wr),
      .wren_b(0),
      .q_a(map_data_out));

  // Renderer
  Renderer renderer(.clk(clk),
                    ._reset(_reset),

                    ._vram_en(_ren_bus_en),
                    ._vram_rd(_ren_bus_rd),
                    ._vram_wr(_ren_bus_wr),
                    ._vram_be(_ren_bus_be),
                    .vram_addr(ren_bus_addr),
                    .vram_data(ren_bus_data),

                    .x(h_pos),
                    .y(v_pos),
                    .vblank(vblank),
                    .hblank(hblank),
                    .rgb_out(ren_rgb_out));

  wire [`REG_DATA_WIDTH * `NUM_MAIN_REGS - 1 : 0] reg_values;

  wire [`REG_DATA_WIDTH-1:0] reg_array [`NUM_MAIN_REGS-1:0];
  genvar i;
  generate
    for (i = 0; i < `NUM_MAIN_REGS; i = i + 1) begin : REGS
      assign reg_array[i] = reg_values[`REG_DATA_WIDTH * (i + 1) - 1:
                                       `REG_DATA_WIDTH * i];
    end
  endgenerate

  // For now, send the values of the register to the lines of the screen, for
  // visual verification.
  // TODO: This test mechanism needs to be changed later.
  assign vga_rgb = (hblank | vblank) ? {`RGB_COLOR_DEPTH {1'b0}}
                                     : {`RGB_COLOR_DEPTH {reg_values[v_pos]}};

  wire main_reg_select = (mpu_addr >= `MAIN_REG_ADDR_BASE) &
                         (mpu_addr < `MAIN_REG_ADDR_BASE + `NUM_MAIN_REGS);
  Registers #(.DATA_WIDTH(`REG_DATA_WIDTH),
              .ADDR_WIDTH(`MAIN_REG_ADDR_WIDTH),
              .NUM_REGS(`NUM_MAIN_REGS))
      registers(.reset(~_reset),
                .en(main_reg_select),
                .rd(~_mpu_rd),
                .wr(~_mpu_wr),
                .be(~_mpu_be),
                .addr(mpu_addr[`MAIN_REG_ADDR_WIDTH-1:0]),
                .data_in(mpu_data),
                .data_out(reg_data_out),
                .values_out(reg_values));

  // VRAM interface logic
  // TODO: the multiplexed VRAM access by both Renderer and MPU here may be too
  // simple.
  wire vram_uses_mpu = ~_mpu_en;
  assign _vram_en = vram_uses_mpu ? _mpu_en : _ren_bus_en;
  assign _vram_wr = vram_uses_mpu ? _mpu_wr : _ren_bus_wr;
  assign _vram_rd = vram_uses_mpu ? _mpu_rd : _ren_bus_rd;
  assign _vram_be = vram_uses_mpu ? _mpu_be : _ren_bus_be;
  assign vram_addr = vram_uses_mpu ? mpu_addr : ren_bus_addr;

  assign vram_data = vram_uses_mpu ? mpu_data : {`VRAM_DATA_WIDTH {1'bz}};
  assign ren_bus_data = vram_data;

endmodule
